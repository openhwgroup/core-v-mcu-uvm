// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_CVMCU_EVENT_FTDECS_SV__
`define __UVMA_CVMCU_EVENT_FTDECS_SV__


typedef class uvma_cvmcu_event_cfg_c     ;
typedef class uvma_cvmcu_event_cntxt_c   ;
typedef class uvma_cvmcu_event_mon_trn_c ;
typedef class uvma_cvmcu_event_seq_item_c;
typedef class uvma_cvmcu_event_phy_mon_trn_c;
typedef class uvma_cvmcu_event_sys_phy_seq_item_c;
typedef class uvma_cvmcu_event_core_phy_seq_item_c;
typedef class uvma_cvmcu_event_mon_vseq_c ;
typedef class uvma_cvmcu_event_idle_vseq_c;
typedef class uvma_cvmcu_event_core_drv_vseq_c;
typedef class uvma_cvmcu_event_sys_drv_vseq_c;


`endif // __UVMA_CVMCU_EVENT_FTDECS_SV__