// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_APB_TIMER_SS_TDEFS_SV__
`define __UVME_APB_TIMER_SS_TDEFS_SV__


// Add tdefs, enums and structs here
// Ex: typedef bit [(`UVME_APB_TIMER_SS_ABC_MAX_WIDTH-1):0]  uvme_apb_timer_ss_abc_b_t;
// Ex: typedef enum {
//        UVME_APB_TIMER_SS_EXAMPLE_ABC
//     } uvme_apb_timer_ss_example_enum;
// Ex: typedef struct {
//        bit [2:0]  abc;
//        logic      xyz;
//     } uvme_apb_timer_ss_example_struct;


`endif // __UVME_APB_TIMER_SS_TDEFS_SV__