// Copyright 2023 Acme Enterprises
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_TCOUNTER_B_MACROS_SVH__
`define __UVMA_TCOUNTER_B_MACROS_SVH__




`endif // __UVMA_TCOUNTER_B_MACROS_SVH__