// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_CVMCU_CPI_ST_FTDECS_SV__
`define __UVME_CVMCU_CPI_ST_FTDECS_SV__


typedef class uvme_cvmcu_cpi_st_cfg_c  ;
typedef class uvme_cvmcu_cpi_st_cntxt_c;


`endif // __UVME_CVMCU_CPI_ST_FTDECS_SV__