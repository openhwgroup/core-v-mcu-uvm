// Copyright 2022 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_CVMCU_INTR_ST_CHKR_SV__
`define __UVME_CVMCU_INTR_ST_CHKR_SV__


/**
 * Encapsulates assertions targeting uvme_cvmcu_intr_st interfaces.
 * This module must be bound to interfaces in a test bench.
 */
module uvme_cvmcu_intr_st_chkr (
      uvma_cvmcu_intr_if  active_if ,
      uvma_cvmcu_intr_if  passive_if
);

   // TODO Add assertions to uvme_cvmcu_intr_st_chkr

endmodule : uvme_cvmcu_intr_st_chkr


`endif // __UVME_CVMCU_INTR_ST_CHKR_SV__
