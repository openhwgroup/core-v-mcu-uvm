// Copyright 2022 Datum Technology Corporation
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
// Licensed under the Solderpad Hardware License v 2.1 (the "License"); you may not use this file except in compliance
// with the License, or, at your option, the Apache License version 2.0.  You may obtain a copy of the License at
//                                        https://solderpad.org/licenses/SHL-2.1/
// Unless required by applicable law or agreed to in writing, any work distributed under the License is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.  See the License for the
// specific language governing permissions and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_CVMCU_DUT_CHKR_SV__
`define __UVMT_CVMCU_DUT_CHKR_SV__


/**
 * Module encapsulating assertions for CORE-V MCU RTL DUT wrapper.  All ports are SV interfaces.
 */
module uvmt_cvmcu_dut_chkr(
   uvma_obi_if  obi_if,
   uvmt_cvmcu_probe_if  probe_if
);
   
   // TODO Add assertions to uvmt_cvmcu_dut_chkr
   
endmodule : uvmt_cvmcu_dut_chkr


`endif // __UVMT_CVMCU_DUT_CHKR_SV__
