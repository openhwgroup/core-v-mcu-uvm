// Copyright 2022 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_UDMA_CTRL_DP_IN_IF_CHKR_SV__
`define __UVMA_UDMA_CTRL_DP_IN_IF_CHKR_SV__


/**
 * Encapsulates assertions targeting uvma_udma_ctrl_dp_in_if.
 * This module must be bound to an interface in a test bench.
 * @ingroup uvma_udma_ctrl_dp_in_misc
 */
module uvma_udma_ctrl_dp_in_if_chkr (
   uvma_udma_ctrl_dp_in_if  udma_ctrl_dp_in_if
);

   // TODO Add assertions to uvma_udma_ctrl_dp_in_if_chkr

endmodule : uvma_udma_ctrl_dp_in_if_chkr


`endif // __UVMA_UDMA_CTRL_DP_IN_IF_CHKR_SV__
