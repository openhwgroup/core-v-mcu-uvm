// Copyright 2022 Datum Technology Corporation
// Copyright 2022 Low Power Futures
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_APB_TIMER_REG_BIT_BASH_VSEQ_IGNORE_LIST_SV__
`define __UVME_APB_TIMER_REG_BIT_BASH_VSEQ_IGNORE_LIST_SV__


string  bb_ignore_list[$] = '{
   // TODO Add registers and/or register blocks to ignore list for automated bit-bash testing
   //      Ex: "reg_name"     , // One register at a time
   //      Ex: "reg_name.abc*", // One register field at a time
   "cfg_reg_hi",
   "cfg_reg_low"
};


`endif // __UVME_APB_TIMER_REG_BIT_BASH_VSEQ_IGNORE_LIST_SV__
