// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_CVMCU_CPI_ST_MACROS_SV__
`define __UVMT_CVMCU_CPI_ST_MACROS_SV__


`ifndef UVMT_CVMCU_CPI_ST_DATA_WIDTH
   `define UVMT_CVMCU_CPI_ST_DATA_WIDTH 12
`endif



`endif // __UVMT_CVMCU_CPI_ST_MACROS_SV__