// Copyright 2022 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_CVMCU_INTR_IF_CHKR_SV__
`define __UVMA_CVMCU_INTR_IF_CHKR_SV__


/**
 * Encapsulates assertions targeting uvma_cvmcu_intr_if.
 * This module must be bound to an interface in a test bench.
 */
module uvma_cvmcu_intr_if_chkr (
   uvma_cvmcu_intr_if  cvmcu_intr_if
);

   // TODO Add assertions to uvma_cvmcu_intr_if_chkr

endmodule : uvma_cvmcu_intr_if_chkr


`endif // __UVMA_CVMCU_INTR_IF_CHKR_SV__
