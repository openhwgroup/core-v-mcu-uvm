// Copyright 2022 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_CVMCU_INTR_ST_CONSTANTS_SV__
`define __UVME_CVMCU_INTR_ST_CONSTANTS_SV__


// Add constants here
// Ex: const int unsigned  uvme_cvmcu_intr_st_my_cons = 10; ///< Describe me!


`endif // __UVME_CVMCU_INTR_ST_CONSTANTS_SV__
