// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_CVMCU_IO_MACROS_SV__
`define __UVMA_CVMCU_IO_MACROS_SV__


`define UVMA_CVMCU_IO_DATA_MIN_SIZE  1
`define UVMA_CVMCU_IO_DATA_MAX_SIZE  `UVM_PACKER_MAX_BYTES


`endif // __UVMA_CVMCU_IO_MACROS_SV__