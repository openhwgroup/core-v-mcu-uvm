// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_CVMCU_CHIP_MACROS_SVH__
`define __UVME_CVMCU_CHIP_MACROS_SVH__


// Add preprocessor macros here
// Ex: `ifndef UVME_CVMCU_CHIP_ABC
//        `define UVME_CVMCU_CHIP_ABC 32
//     `endif


`endif // __UVME_CVMCU_CHIP_MACROS_SVH__