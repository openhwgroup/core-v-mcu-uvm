// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_TPRESCALER_B_TDEFS_SV__
`define __UVMA_TPRESCALER_B_TDEFS_SV__



/// @name Logic vectors
/// @{
typedef logic [31:0]  uvma_tprescaler_b_compare_value_i_l_t; ///<  logic vector
typedef logic [31:0]  uvma_tprescaler_b_counter_value_i_l_t; ///<  logic vector
typedef logic [31:0]  uvma_tprescaler_b_counter_value_o_l_t; ///<  logic vector
/// @}

/// @name Bit vectors
/// @{
typedef bit [31:0]  uvma_tprescaler_b_compare_value_i_b_t; ///<  bit vector
typedef bit [31:0]  uvma_tprescaler_b_counter_value_i_b_t; ///<  bit vector
typedef bit [31:0]  uvma_tprescaler_b_counter_value_o_b_t; ///<  bit vector
/// @}


`endif // __UVMA_TPRESCALER_B_TDEFS_SV__