// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_CVMCU_CPI_CONSTANTS_SV__
`define __UVMA_CVMCU_CPI_CONSTANTS_SV__


`endif // __UVMA_CVMCU_CPI_CONSTANTS_SV__