// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_CVMCU_CPI_MACROS_SV__
`define __UVMA_CVMCU_CPI_MACROS_SV__


`define UVMA_CVMCU_CPI_DATA_MIN_SIZE  8
`define UVMA_CVMCU_CPI_DATA_MAX_SIZE  1_024
`define UVMA_CVMCU_CPI_DATA_MIN_WIDTH  12
`define UVMA_CVMCU_CPI_DATA_MAX_WIDTH  20


`endif // __UVMA_CVMCU_CPI_MACROS_SV__