// Copyright 2022 Datum Technology Corporation
// Copyright 2022 Low Power Futures
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_APB_TIMER_REG_BIT_BASH_VSEQ_IGNORE_LIST_SV__
`define __UVME_APB_TIMER_REG_BIT_BASH_VSEQ_IGNORE_LIST_SV__


string  bb_ignore_list[$] = '{
   "cfg_reg_hi" ,
   "cfg_reg_low"
};


`endif // __UVME_APB_TIMER_REG_BIT_BASH_VSEQ_IGNORE_LIST_SV__
