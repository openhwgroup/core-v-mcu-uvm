// Copyright 2023 Acme Enterprises
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_TPRESCALER_B_TDEFS_SV__
`define __UVMT_TPRESCALER_B_TDEFS_SV__


// Add enums and structs here
// Ex: typedef bit [(`UVMT_TPRESCALER_B_ABC_MAX_WIDTH-1):0]  uvmt_tprescaler_b_abc_b_t; ///< Describe me!
// Ex: /*
//      * Describe me!
//      */
//     typedef enum {
//        UVMT_TPRESCALER_B_EX_ABC
//     } uvmt_tprescaler_b_ex_enum;
// Ex: /*
//      * Describe me!
//      */
//     typedef struct {
//        bit [2:0]  abc;
//        logic      xyz;
//     } uvmt_tprescaler_b_ex_struct;


`endif // __UVMT_TPRESCALER_B_TDEFS_SV__