// Copyright 2023 Acme Enterprises
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_CVMCU_DBG_SYS_PHY_DRV_SV__
`define __UVMA_CVMCU_DBG_SYS_PHY_DRV_SV__


/**
 * Driver driving CORE-V-MCU Debug Interface Virtual Interface (uvma_cvmcu_dbg_if) SYS PHY.
 * @ingroup uvma_cvmcu_dbg_comps
 */
class uvma_cvmcu_dbg_sys_phy_drv_c extends uvmx_mp_drv_c #(
   .T_MP      (virtual uvma_cvmcu_dbg_if.sys_phy_drv_mp),
   .T_CFG     (uvma_cvmcu_dbg_cfg_c  ),
   .T_CNTXT   (uvma_cvmcu_dbg_cntxt_c),
   .T_SEQ_ITEM(uvma_cvmcu_dbg_sys_phy_seq_item_c)
);

   `uvm_component_utils(uvma_cvmcu_dbg_sys_phy_drv_c)
   `uvmx_mp_drv(sys_phy_drv_mp, sys_phy_drv_cb)

   /**
    * Default constructor.
    */
   function new(string name="uvma_cvmcu_dbg_sys_phy_drv", uvm_component parent=null);
      super.new(name, parent);
   endfunction


   /**
    * Drives SYS PHY Driver clocking block (sys_phy_drv_cb) on each clock cycle.
    */
   virtual task drive_item(ref uvma_cvmcu_dbg_sys_phy_seq_item_c item);
      mp.sys_phy_drv_cb.debug_req_i <= item.debug_req_i;
   endtask

   /**
    * Samples SYS PHY Driver clocking block (sys_phy_drv_cb) after each clock cycle.
    */
   virtual task sample_post_clk(ref uvma_cvmcu_dbg_sys_phy_seq_item_c item);
      item.stoptimer_o = mp.sys_phy_drv_cb.stoptimer_o;
   endtask

endclass : uvma_cvmcu_dbg_sys_phy_drv_c


`endif // __UVMA_CVMCU_DBG_SYS_PHY_DRV_SV__