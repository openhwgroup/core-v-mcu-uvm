// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_TCOUNTER_B_MACROS_SVH__
`define __UVMT_TCOUNTER_B_MACROS_SVH__


// Add preprocessor macros here
// Ex: `ifndef UVMT_TCOUNTER_B_ABC_WIDTH
//        `define UVMT_TCOUNTER_B_ABC_WIDTH 32
//     `endif


`endif // __UVMT_TCOUNTER_B_MACROS_SVH__