// Copyright 2022-2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_CVMCU_TDEFS_SV__
`define __UVMT_CVMCU_TDEFS_SV__


// Add enums and structs here
// Ex: typedef bit [(`UVMT_CVMCU_ABC_MAX_WIDTH-1):0]  uvmt_cvmcu_abc_b_t;
// Ex: typedef enum {
//        UVMT_CVMCU_MY_ABC
//     } uvmt_cvmcu_my_enum;
// Ex: typedef struct {
//        bit [2:0]  abc;
//        logic      xyz;
//     } uvmt_cvmcu_my_struct;


`endif // __UVMT_CVMCU_TDEFS_SV__