// Copyright 2023 Acme Enterprises
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_ADV_TIMER_B_CONSTANTS_SV__
`define __UVME_ADV_TIMER_B_CONSTANTS_SV__


const int unsigned  uvme_adv_timer_b_default_num_items_cons = 10; ///< Default number of Sequence Items to be generated in a Sequence.


`endif // __UVME_ADV_TIMER_B_CONSTANTS_SV__