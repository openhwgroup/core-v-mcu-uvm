// Copyright 2023 Acme Enterprises
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_CVMCU_DBG_ST_CONSTANTS_SV__
`define __UVME_CVMCU_DBG_ST_CONSTANTS_SV__



const int unsigned  uvme_cvmcu_dbg_st_rand_stim_vseq_default_num_items      = 10; ///< Default number of Sequence Items generated by sequences.
const int unsigned  uvme_cvmcu_dbg_st_rand_stim_vseq_default_min_size       =  8; ///< Default minimum packet size for sequences.
const int unsigned  uvme_cvmcu_dbg_st_rand_stim_vseq_default_max_size       = 64; ///< Default maximum packet size for sequences.
const int unsigned  uvme_cvmcu_dbg_st_rand_stim_vseq_default_min_gap        =  0; ///< Default minimum gap for sequences.
const int unsigned  uvme_cvmcu_dbg_st_rand_stim_vseq_default_max_gap        = 10; ///< Default maximum gap for sequences.
const int unsigned  uvme_cvmcu_dbg_st_rand_ill_stim_vseq_default_num_items  = 10; ///< Default number of Sequence Items generated by error sequences.
const int unsigned  uvme_cvmcu_dbg_st_rand_ill_stim_vseq_default_num_errors =  1; ///< Default number of illegal sequence items generated by error sequences.
const int unsigned  uvme_cvmcu_dbg_st_rand_ill_stim_vseq_default_min_size   =  8; ///< Default minimum packet size for error sequences.
const int unsigned  uvme_cvmcu_dbg_st_rand_ill_stim_vseq_default_max_size   = 64; ///< Default maximum packet size for error sequences.
const int unsigned  uvme_cvmcu_dbg_st_rand_ill_stim_vseq_default_min_gap    =  0; ///< Default minimum gap for error sequences.
const int unsigned  uvme_cvmcu_dbg_st_rand_ill_stim_vseq_default_max_gap    = 10; ///< Default maximum gap for error sequences.



`endif // __UVME_CVMCU_DBG_ST_CONSTANTS_SV__