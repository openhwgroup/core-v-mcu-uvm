// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_TCOUNTER_B_CONSTANTS_SV__
`define __UVME_TCOUNTER_B_CONSTANTS_SV__


`endif // __UVME_TCOUNTER_B_CONSTANTS_SV__