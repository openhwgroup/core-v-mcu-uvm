// Copyright 2022 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_UDMA_TX_DP_IN_MACROS_SVH__
`define __UVMA_UDMA_TX_DP_IN_MACROS_SVH__


// Add preprocessor macros here
// Ex: `ifndef UVMA_UDMA_TX_DP_IN_ABC_MAX_WIDTH
//        `define UVMA_UDMA_TX_DP_IN_ABC_MAX_WIDTH 32
//     `endif


`endif // __UVMA_UDMA_TX_DP_IN_MACROS_SVH__
