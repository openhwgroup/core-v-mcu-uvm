// Copyright 2023 Acme Enterprises
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_CVMCU_IO_IF_CHKR_SV__
`define __UVMA_CVMCU_IO_IF_CHKR_SV__


/**
 * Encapsulates assertions targeting uvma_cvmcu_io_if.
 * @ingroup uvma_cvmcu_io_misc
 */
module uvma_cvmcu_io_if_chkr(
   uvma_cvmcu_io_if  cvmcu_io_if  ///< Target interface handle
);

   // TODO Add assertions to uvma_cvmcu_io_if_chkr

endmodule : uvma_cvmcu_io_if_chkr


`endif // __UVMA_CVMCU_IO_IF_CHKR_SV__