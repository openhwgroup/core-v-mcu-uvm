// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_TPRESCALER_B_FTDECS_SV__
`define __UVME_TPRESCALER_B_FTDECS_SV__


`endif // __UVME_TPRESCALER_B_FTDECS_SV__