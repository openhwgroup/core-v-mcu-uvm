// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_CVMCU_DBG_IF_CHKR_SV__
`define __UVMA_CVMCU_DBG_IF_CHKR_SV__


/**
 * Encapsulates assertions targeting uvma_cvmcu_dbg_if.
 * @ingroup uvma_cvmcu_dbg_misc
 */
module uvma_cvmcu_dbg_if_chkr(
   uvma_cvmcu_dbg_if  cvmcu_dbg_if  ///< Target interface handle
);

   // TODO Add assertions to uvma_cvmcu_dbg_if_chkr

endmodule : uvma_cvmcu_dbg_if_chkr


`endif // __UVMA_CVMCU_DBG_IF_CHKR_SV__