// Copyright 2022 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_UDMA_RX_TDEFS_SV__
`define __UVMT_UDMA_RX_TDEFS_SV__


// Add tdefs, enums and structs here
// Ex: typedef bit [(`UVMT_UDMA_RX_ABC_MAX_WIDTH-1):0]  uvmt_udma_rx_abc_b_t;
// Ex: typedef enum {
//        UVMT_UDMA_RX_MY_ABC
//     } uvmt_udma_rx_my_enum;
// Ex: typedef struct {
//        bit [2:0]  abc;
//        logic      xyz;
//     } uvmt_udma_rx_my_struct;


`endif // __UVMT_UDMA_RX_TDEFS_SV__
