// Copyright 2023 Acme Enterprises
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_CVMCU_CHIP_TDEFS_SV__
`define __UVMT_CVMCU_CHIP_TDEFS_SV__


// Add enums and structs here
// Ex: typedef bit [(`UVMT_CVMCU_CHIP_ABC_MAX_WIDTH-1):0]  uvmt_cvmcu_chip_abc_b_t;
// Ex: typedef enum {
//        UVMT_CVMCU_CHIP_EXAMPLE_ABC
//     } uvmt_cvmcu_chip_example_enum;
// Ex: typedef struct {
//        bit [2:0]  abc;
//        logic      xyz;
//     } uvmt_cvmcu_chip_example_struct;


`endif // __UVMT_CVMCU_CHIP_TDEFS_SV__