// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_CVMCU_CHIP_FTDECS_SV__
`define __UVME_CVMCU_CHIP_FTDECS_SV__



`endif // __UVME_CVMCU_CHIP_FTDECS_SV__