// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_TCOUNTER_B_FTDECS_SV__
`define __UVMA_TCOUNTER_B_FTDECS_SV__


typedef class uvma_tcounter_b_cfg_c         ;
typedef class uvma_tcounter_b_cntxt_c       ;
typedef class uvma_tcounter_b_seq_item_c    ;
typedef class uvma_tcounter_b_cp_seq_item_c ;
typedef class uvma_tcounter_b_dpi_seq_item_c;
typedef class uvma_tcounter_b_dpo_seq_item_c;
typedef class uvma_tcounter_b_mon_seq_c     ;
typedef class uvma_tcounter_b_idle_seq_c    ;
typedef class uvma_tcounter_b_in_drv_seq_c  ;
typedef class uvma_tcounter_b_out_drv_seq_c ;


`endif // __UVMA_TCOUNTER_B_FTDECS_SV__