// Copyright 2022 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_CVMCU_INTR_ST_MACROS_SV__
`define __UVMT_CVMCU_INTR_ST_MACROS_SV__


// Add preprocessor macros here
// Ex: `ifndef UVMT_CVMCU_INTR_ST_ABC_MAX_WIDTH
//        `define UVMT_CVMCU_INTR_ST_ABC_MAX_WIDTH 32
//     `endif


`endif // __UVMT_CVMCU_INTR_ST_MACROS_SV__
