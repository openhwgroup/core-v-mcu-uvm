// Copyright 2022-2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_APB_TIMER_TDEFS_SV__
`define __UVMT_APB_TIMER_TDEFS_SV__


// Add enums and structs here
// Ex: typedef bit [(`UVMT_APB_TIMER_ABC_MAX_WIDTH-1):0]  uvmt_apb_timer_abc_b_t;
// Ex: typedef enum {
//        UVMT_APB_TIMER_MY_ABC
//     } uvmt_apb_timer_my_enum;
// Ex: typedef struct {
//        bit [2:0]  abc;
//        logic      xyz;
//     } uvmt_apb_timer_my_struct;


`endif // __UVMT_APB_TIMER_TDEFS_SV__