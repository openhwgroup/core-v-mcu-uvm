// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_APB_TIMER_SS_MACROS_SVH__
`define __UVME_APB_TIMER_SS_MACROS_SVH__


// Add preprocessor macros here
// Ex: `ifndef UVME_APB_TIMER_SS_ABC
//        `define UVME_APB_TIMER_SS_ABC 32
//     `endif


`endif // __UVME_APB_TIMER_SS_MACROS_SVH__