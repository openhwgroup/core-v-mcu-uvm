// Copyright 2023 Acme Enterprises
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_CVMCU_CPI_ST_TDEFS_SV__
`define __UVMT_CVMCU_CPI_ST_TDEFS_SV__


// Add enums and structs here
// Ex: typedef bit [(`UVMT__ST_ABC_MAX_WIDTH-1):0]  uvmt_cvmcu_cpi_st_abc_b_t; ///< Describe me!
// Ex: /*
//      * Describe me!
//      */
//     typedef enum {
//        UVMT__ST_EX_ABC
//     } uvmt_cvmcu_cpi_st_ex_enum;
// Ex: /*
//      * Describe me!
//      */
//     typedef struct {
//        bit [2:0]  abc;
//        logic      xyz;
//     } uvmt_cvmcu_cpi_st_ex_struct;


`endif // __UVMT_CVMCU_CPI_ST_TDEFS_SV__