// Copyright 2023 Acme Enterprises
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_CVMCU_DBG_ST_MACROS_SV__
`define __UVMT_CVMCU_DBG_ST_MACROS_SV__


// Add preprocessor macros here
// Ex: `ifndef UVMT_CVMCU_DBG_ST_ABC_WIDTH
//        `define UVMT_CVMCU_DBG_ST_ABC_WIDTH 32
//     `endif



`endif // __UVMT_CVMCU_DBG_ST_MACROS_SV__