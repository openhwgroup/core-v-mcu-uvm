// Copyright 2023 Acme Enterprises
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_TPRESCALER_B_CONSTANTS_SV__
`define __UVME_TPRESCALER_B_CONSTANTS_SV__


const int unsigned  uvme_tprescaler_b_default_num_items_cons = 10; ///< Default number of Sequence Items to be generated in a Sequence.


`endif // __UVME_TPRESCALER_B_CONSTANTS_SV__