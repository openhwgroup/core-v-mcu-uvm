// Copyright 2023 Acme Enterprises
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_TCOUNTER_B_CONSTANTS_SV__
`define __UVMA_TCOUNTER_B_CONSTANTS_SV__




`endif // __UVMA_TCOUNTER_B_CONSTANTS_SV__