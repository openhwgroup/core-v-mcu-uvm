// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_CVMCU_CHIP_TDEFS_SV__
`define __UVME_CVMCU_CHIP_TDEFS_SV__



`endif // __UVME_CVMCU_CHIP_TDEFS_SV__