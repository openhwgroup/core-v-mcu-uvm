// Copyright 2022 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_UDMA_RX_CONSTANTS_SV__
`define __UVME_UDMA_RX_CONSTANTS_SV__


const int unsigned  uvme_udma_rx_default_clk_frequency = 100_000_000; ///< Clock agent frequency (Hz)


`endif // __UVME_UDMA_RX_CONSTANTS_SV__
