// Copyright 2023 Acme Enterprises
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_TPRESCALER_B_CONSTANTS_SV__
`define __UVMA_TPRESCALER_B_CONSTANTS_SV__




`endif // __UVMA_TPRESCALER_B_CONSTANTS_SV__