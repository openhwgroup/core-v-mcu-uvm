// Copyright 2022 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_CVMCU_MACROS_SVH__
`define __UVMT_CVMCU_MACROS_SVH__


// Add preprocessor macros here
// Ex: `ifndef UVMT_CVMCU_ABC_MAX_WIDTH
//        `define UVMT_CVMCU_ABC_MAX_WIDTH 32
//     `endif


`endif // __UVMT_CVMCU_MACROS_SVH__