// Copyright 2022 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_CVMCU_INTR_CONSTANTS_SV__
`define __UVMA_CVMCU_INTR_CONSTANTS_SV__


// Add constants here
// Ex: const int unsigned  uvma_cvmcu_intr_my_cons = 10;


`endif // __UVMA_CVMCU_INTR_CONSTANTS_SV__
