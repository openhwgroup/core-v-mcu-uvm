// Copyright 2024 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_APB_ADV_TIMER_SS_BASE_TEST_WORKAROUNDS_SV__
`define __UVMT_APB_ADV_TIMER_SS_BASE_TEST_WORKAROUNDS_SV__


// Temporary configuration constraints here (this file should be empty by the end of the project).


`endif // __UVMT_APB_ADV_TIMER_SS_BASE_TEST_WORKAROUNDS_SV__