// Copyright 2022 Datum Technology Corporation
// Copyright 2022 Low Power Futures
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_APB_ADV_TIMER_REG_HW_RESET_VSEQ_IGNORE_LIST_SV__
`define __UVME_APB_ADV_TIMER_REG_HW_RESET_VSEQ_IGNORE_LIST_SV__


string  ignore_list[$] = '{
   // TODO Add registers and/or register blocks to ignore list for automated testing of reset values
   //      Ex: "block_name.reg_name", // One register at a time
   //      Ex: "block_name.*", // One block at a time
};


`endif // __UVME_APB_ADV_TIMER_REG_HW_RESET_VSEQ_IGNORE_LIST_SV__
