// Copyright 2022 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_CVMCU_INTR_ST_DUT_CHKR_SV__
`define __UVMT_CVMCU_INTR_ST_DUT_CHKR_SV__


/**
 * Module encapsulating assertions for the CORE-V MCU Interrupt UVM Agent Self-Test DUT wrapper (uvmt_cvmcu_intr_st_dut_wrap).
 */
module uvmt_cvmcu_intr_st_dut_chkr (
   uvma_cvmcu_intr_if  active_if , ///< Active agent interface
   uvma_cvmcu_intr_if  passive_if ///< Passive agent interface
);

   // TODO Add assertions to uvmt_cvmcu_intr_st_dut_chkr

endmodule : uvmt_cvmcu_intr_st_dut_chkr


`endif // __UVMT_CVMCU_INTR_ST_DUT_CHKR_SV__
