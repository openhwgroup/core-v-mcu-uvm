// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_TCOUNTER_B_FTDECS_SV__
`define __UVMT_TCOUNTER_B_FTDECS_SV__


`endif // __UVMT_TCOUNTER_B_FTDECS_SV__