// Copyright 2022-2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_APB_ADV_TIMER_CONSTANTS_SV__
`define __UVME_APB_ADV_TIMER_CONSTANTS_SV__


const longint unsigned  uvme_apb_adv_timer_default_reg_block_base_address = 64'h0000_0000_0000_0000; ///< Register block base address
const int unsigned      uvme_apb_adv_timer_reg_block_reg_n_bytes          = 4; ///< Width of registers (bytes)


`endif // __UVME_APB_ADV_TIMER_CONSTANTS_SV__