// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_ADV_TIMER_B_MACROS_SVH__
`define __UVMT_ADV_TIMER_B_MACROS_SVH__


`ifndef UVMT_ADV_TIMER_B_NUM_BITS
   `define UVMT_ADV_TIMER_B_NUM_BITS 16
`endif
`ifndef UVMT_ADV_TIMER_B_N_EXTSIG
   `define UVMT_ADV_TIMER_B_N_EXTSIG 32
`endif


`endif // __UVMT_ADV_TIMER_B_MACROS_SVH__