// Copyright 2023 Acme Enterprises
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_APB_ADV_TIMER_SS_REG_IGNORE_LISTS_SV__
`define __UVME_APB_ADV_TIMER_SS_REG_IGNORE_LISTS_SV__


string  uvme_apb_adv_timer_ss_all_reg_mem_ignore_list[$] = '{
};

string  uvme_apb_adv_timer_ss_reg_hw_reset_ignore_list[$] = '{
};

string  uvme_apb_adv_timer_ss_reg_bit_bash_ignore_list[$] = '{
};

string  uvme_apb_adv_timer_ss_reg_access_ignore_list[$] = '{
};

string  uvme_apb_adv_timer_ss_mem_access_ignore_list[$] = '{
};

string  uvme_apb_adv_timer_ss_shared_access_ignore_list[$] = '{
};

string  uvme_apb_adv_timer_ss_mem_walk_access_ignore_list[$] = '{
};


`endif // __UVME_APB_ADV_TIMER_SS_REG_IGNORE_LISTS_SV__