// Copyright 2022 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_CVMCU_INTR_ST_TDEFS_SV__
`define __UVMT_CVMCU_INTR_ST_TDEFS_SV__


// Add enums and structs here
// Ex: typedef enum {
//        UVMT_CVMCU_INTR_ST_MY_ABC
//     } uvmt_cvmcu_intr_st_my_enum;
// Ex: typedef struct {
//        bit [2:0]  abc;
//        logic      xyz;
//     } uvmt_cvmcu_intr_st_my_struct;


`endif // __UVMT_CVMCU_INTR_ST_TDEFS_SV__
