// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_TCOUNTER_B_DPI_DRV_SV__
`define __UVMA_TCOUNTER_B_DPI_DRV_SV__


/**
 * Driver driving uvma_tcounter_b_if with Data Plane Input Sequence Items (uvma_tcounter_b_dpi_seq_item_c).
 * @ingroup uvma_tcounter_b_comps
 */
class uvma_tcounter_b_dpi_drv_c extends uvmx_mp_drv_c #(
   .T_MP      (virtual uvma_tcounter_b_if.dpi_drv_mp),
   .T_CFG     (uvma_tcounter_b_cfg_c                ),
   .T_CNTXT   (uvma_tcounter_b_cntxt_c              ),
   .T_SEQ_ITEM(uvma_tcounter_b_dpi_seq_item_c       )
);

   `uvm_component_utils(uvma_tcounter_b_dpi_drv_c)
   `uvmx_mp_drv(dpi_drv_mp, dpi_drv_cb)


   /**
    * Default constructor.
    */
   function new(string name="uvma_tcounter_b_dpi_drv", uvm_component parent=null);
      super.new(name, parent);
   endfunction

   /**
    * Drives the Data Plane Input driver clocking block (dpi_drv_cb) on each clock cycle.
    */
   virtual task drive_item(ref uvma_tcounter_b_dpi_seq_item_c item);
      `uvmx_mp_drv_signal(item, write_counter_i)
      `uvmx_mp_drv_signal(item, counter_value_i)
   endtask


endclass : uvma_tcounter_b_dpi_drv_c


`endif // __UVMA_TCOUNTER_B_DPI_DRV_SV__