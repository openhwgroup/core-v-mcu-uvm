// Copyright 2022-2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_CVMCU_TDEFS_SV__
`define __UVME_CVMCU_TDEFS_SV__


// TODO Add scoreboard specialization(s)
//      Ex: typedef uvml_sb_simplex_c#(
//             .T_CNTXT(uvme_cvmcu_sb_cntxt_c),
//             .T_TRN  (uvma_cvmcu_mon_trn_c )
//          ) uvme_cvmcu_sb_simplex_c;

// Add tdefs, enums and structs here
// Ex: typedef bit [(`UVME_CVMCU_ABC_MAX_WIDTH-1):0]  uvme_cvmcu_abc_b_t;
// Ex: typedef enum {
//        UVME_CVMCU_MY_ABC
//     } uvme_cvmcu_my_enum;
// Ex: typedef struct {
//        bit [2:0]  abc;
//        logic      xyz;
//     } uvme_cvmcu_my_struct;


`endif // __UVME_CVMCU_TDEFS_SV__