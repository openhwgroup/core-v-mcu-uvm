// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_CVMCU_EVENT_IF_CHKR_SV__
`define __UVMA_CVMCU_EVENT_IF_CHKR_SV__


/**
 * Encapsulates assertions targeting uvma_cvmcu_event_if.
 * @ingroup uvma_cvmcu_event_misc
 */
module uvma_cvmcu_event_if_chkr(
   uvma_cvmcu_event_if  cvmcu_event_if  ///< Target interface handle
);

   // TODO Add assertions and/or functional coverage to uvma_cvmcu_event_if_chkr

endmodule : uvma_cvmcu_event_if_chkr


`endif // __UVMA_CVMCU_EVENT_IF_CHKR_SV__