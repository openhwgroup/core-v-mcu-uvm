// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_ADV_TIMER_B_MACROS_SVH__
`define __UVME_ADV_TIMER_B_MACROS_SVH__


// Add preprocessor macros here
// Ex: `ifndef UVME_ADV_TIMER_B_ABC
//        `define UVME_ADV_TIMER_B_ABC 32
//     `endif


`endif // __UVME_ADV_TIMER_B_MACROS_SVH__