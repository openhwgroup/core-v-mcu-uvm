// Copyright 2022 Datum Technology Corporation
// Copyright 2022 Low Power Futures
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_APB_TIMER_MACROS_SVH__
`define __UVME_APB_TIMER_MACROS_SVH__


// Add preprocessor macros here
// Ex: `ifndef UVME_APB_TIMER_ABC
//        `define UVME_APB_TIMER_ABC 32
//     `endif


`endif // __UVME_APB_TIMER_MACROS_SVH__
