// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_CVMCU_CHIP_MACROS_SVH__
`define __UVMT_CVMCU_CHIP_MACROS_SVH__


`ifndef UVMT_CVMCU_CHIP_USE_CORES
   `define UVMT_CVMCU_CHIP_USE_CORES 0
`endif



`endif // __UVMT_CVMCU_CHIP_MACROS_SVH__