// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_CVMCU_CHIP_FTDECS_SV__
`define __UVME_CVMCU_CHIP_FTDECS_SV__


typedef class uvme_cvmcu_chip_udma_uart_seq_c;


`endif // __UVME_CVMCU_CHIP_FTDECS_SV__
