// Copyright 2023 Acme Enterprises
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_ADV_TIMER_B_IF_CHKR_SV__
`define __UVMA_ADV_TIMER_B_IF_CHKR_SV__


/**
 * Module encapsulating assertions targeting  Block Agent interface.
 * @ingroup uvma_adv_timer_b_pkg
 */
module uvma_adv_timer_b_if_chkr (
   uvma_adv_timer_b_if  agent_if ///< Target interface
);

   // TODO Add assertions to uvme_adv_timer_b_chkr

endmodule : uvma_adv_timer_b_if_chkr


`endif // __UVMA_ADV_TIMER_B_IF_CHKR_SV__