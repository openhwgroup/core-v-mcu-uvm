// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_TPRESCALER_B_IF_CHKR_SV__
`define __UVMA_TPRESCALER_B_IF_CHKR_SV__


/**
 * Module encapsulating assertions targeting Timer unit prescaler Block Agent interface.
 * @ingroup uvma_tprescaler_b_pkg
 */
module uvma_tprescaler_b_if_chkr (
   uvma_tprescaler_b_if  agent_if ///< Target interface
);

   // TODO Add assertions and/or functional coverage to uvme_tprescaler_b_chkr

endmodule


`endif // __UVMA_TPRESCALER_B_IF_CHKR_SV__