// Copyright 2022 Datum Technology Corporation
// Copyright 2022 Low Power Futures
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_APB_TIMER_MACROS_SVH__
`define __UVMT_APB_TIMER_MACROS_SVH__


// Add preprocessor macros here
// Ex: `ifndef UVMT_APB_TIMER_ABC_MAX_WIDTH
//        `define UVMT_APB_TIMER_ABC_MAX_WIDTH 32
//     `endif


`endif // __UVMT_APB_TIMER_MACROS_SVH__
