// Copyright 2023 Acme Enterprises
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_CVMCU_DBG_ST_MACROS_SV__
`define __UVME_CVMCU_DBG_ST_MACROS_SV__


// Add preprocessor macros here
// Ex: `ifndef UVME__ST_ABC
//        `define UVME__ST_ABC 32
//     `endif


`endif // __UVME_CVMCU_DBG_ST_MACROS_SV__