// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_TCOUNTER_B_CONSTANTS_SV__
`define __UVME_TCOUNTER_B_CONSTANTS_SV__


const int unsigned  uvme_tcounter_b_default_num_items_cons = 10; ///< Default number of Sequence Items to be generated in a Sequence.


`endif // __UVME_TCOUNTER_B_CONSTANTS_SV__