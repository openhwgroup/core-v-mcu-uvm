// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_CVMCU_CHIP_TDEFS_SV__
`define __UVME_CVMCU_CHIP_TDEFS_SV__


// Add tdefs, enums and structs here
// Ex: typedef bit [(`UVME_CVMCU_CHIP_ABC_MAX_WIDTH-1):0]  uvme_cvmcu_chip_abc_b_t;
// Ex: typedef enum {
//        UVME_CVMCU_CHIP_EXAMPLE_ABC
//     } uvme_cvmcu_chip_example_enum;
// Ex: typedef struct {
//        bit [2:0]  abc;
//        logic      xyz;
//     } uvme_cvmcu_chip_example_struct;


`endif // __UVME_CVMCU_CHIP_TDEFS_SV__