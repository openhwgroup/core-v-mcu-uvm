// Copyright 2023 Acme Enterprises
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_CVMCU_IO_MACROS_SV__
`define __UVMA_CVMCU_IO_MACROS_SV__


`define UVMA_CVMCU_IO_DATA_MIN_SIZE  8
`define UVMA_CVMCU_IO_DATA_MAX_SIZE  1_024


`endif // __UVMA_CVMCU_IO_MACROS_SV__