// Copyright 2022 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_CVMCU_INTR_TDEFS_SV__
`define __UVMA_CVMCU_INTR_TDEFS_SV__


// Add enums and structs here
// Ex: typedef bit [(`UVMA_CVMCU_INTR_ABC_MAX_WIDTH-1):0]  uvma_cvmcu_intr_abc_b_t;
// Ex: typedef enum {
//        UVMA_CVMCU_INTR_MY_ABC
//     } uvma_cvmcu_intr_my_enum;
// Ex: typedef struct {
//        bit [2:0]  abc;
//        logic      xyz;
//     } uvma_cvmcu_intr_my_struct;


`endif // __UVMA_CVMCU_INTR_TDEFS_SV__
