// Copyright 2023 Acme Enterprises
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_ADV_TIMER_B_MACROS_SVH__
`define __UVMA_ADV_TIMER_B_MACROS_SVH__


`define UVMA_ADV_TIMER_B_NUM_BITS_MIN  16
`define UVMA_ADV_TIMER_B_NUM_BITS_MAX  64
`define UVMA_ADV_TIMER_B_N_EXTSIG_MIN  32
`define UVMA_ADV_TIMER_B_N_EXTSIG_MAX  64


`endif // __UVMA_ADV_TIMER_B_MACROS_SVH__