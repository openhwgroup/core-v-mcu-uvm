// Copyright 2022-2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_CVMCU_CONSTANTS_SV__
`define __UVME_CVMCU_CONSTANTS_SV__


const longint unsigned  uvme_cvmcu_default_reg_block_base_address = `UVM_REG_ADDR_WIDTH'h0000_0000; ///< Register block base address
const int unsigned      uvme_cvmcu_reg_block_reg_n_bytes          = 4; ///< Width of registers (bytes)


`endif // __UVME_CVMCU_CONSTANTS_SV__
