// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_APB_TIMER_SS_TDEFS_SV__
`define __UVMT_APB_TIMER_SS_TDEFS_SV__


// Add enums and structs here
// Ex: typedef bit [(`UVMT_APB_TIMER_SS_ABC_MAX_WIDTH-1):0]  uvmt_apb_timer_ss_abc_b_t;
// Ex: typedef enum {
//        UVMT_APB_TIMER_SS_EXAMPLE_ABC
//     } uvmt_apb_timer_ss_example_enum;
// Ex: typedef struct {
//        bit [2:0]  abc;
//        logic      xyz;
//     } uvmt_apb_timer_ss_example_struct;


`endif // __UVMT_APB_TIMER_SS_TDEFS_SV__