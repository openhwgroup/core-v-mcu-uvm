// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_CVMCU_CPI_FTDECS_SV__
`define __UVMA_CVMCU_CPI_FTDECS_SV__


typedef class uvma_cvmcu_cpi_cfg_c     ;
typedef class uvma_cvmcu_cpi_cntxt_c   ;
typedef class uvma_cvmcu_cpi_mon_trn_c ;
typedef class uvma_cvmcu_cpi_seq_item_c;
typedef class uvma_cvmcu_cpi_phy_mon_trn_c;
typedef class uvma_cvmcu_cpi_tx_phy_seq_item_c;
typedef class uvma_cvmcu_cpi_rx_phy_seq_item_c;
typedef class uvma_cvmcu_cpi_mon_vseq_c ;
typedef class uvma_cvmcu_cpi_idle_vseq_c;
typedef class uvma_cvmcu_cpi_tx_drv_vseq_c;
typedef class uvma_cvmcu_cpi_rx_drv_vseq_c;


`endif // __UVMA_CVMCU_CPI_FTDECS_SV__