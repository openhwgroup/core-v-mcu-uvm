// Copyright 2023 Acme Enterprises
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_TCOUNTER_B_MACROS_SVH__
`define __UVME_TCOUNTER_B_MACROS_SVH__


// Add preprocessor macros here
// Ex: `ifndef UVME_TCOUNTER_B_ABC
//        `define UVME_TCOUNTER_B_ABC 32
//     `endif


`endif // __UVME_TCOUNTER_B_MACROS_SVH__