// Copyright 2024 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_APB_ADV_TIMER_SS_FTDECS_SV__
`define __UVME_APB_ADV_TIMER_SS_FTDECS_SV__


typedef class uvme_apb_adv_timer_ss_reset_seq_c;
typedef class uvme_apb_adv_timer_ss_cfg_seq_c;



`endif // __UVME_APB_ADV_TIMER_SS_FTDECS_SV__