// Copyright 2022 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_UDMA_CTRL_DP_IN_CONSTANTS_SV__
`define __UVMA_UDMA_CTRL_DP_IN_CONSTANTS_SV__


// Add constants here
// Ex: const int unsigned  uvma_udma_ctrl_dp_in_my_cons = 10;


`endif // __UVMA_UDMA_CTRL_DP_IN_CONSTANTS_SV__
