// Copyright 2024 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_APB_TIMER_SS_MACROS_SVH__
`define __UVMT_APB_TIMER_SS_MACROS_SVH__


// Add preprocessor macros here
// Ex: `ifndef UVMT_APB_TIMER_SS_ABC_WIDTH
//        `define UVMT_APB_TIMER_SS_ABC_WIDTH 32
//     `endif



`endif // __UVMT_APB_TIMER_SS_MACROS_SVH__