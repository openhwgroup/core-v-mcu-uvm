// Copyright 2022 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_UDMA_TX_MACROS_SVH__
`define __UVMT_UDMA_TX_MACROS_SVH__


// Add preprocessor macros here
// Ex: `ifndef UVMT_UDMA_TX_ABC_MAX_WIDTH
//        `define UVMT_UDMA_TX_ABC_MAX_WIDTH 32
//     `endif


`endif // __UVMT_UDMA_TX_MACROS_SVH__
