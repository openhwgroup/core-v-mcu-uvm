// Copyright 2022-2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_APB_TIMER_TDEFS_SV__
`define __UVME_APB_TIMER_TDEFS_SV__


// TODO Add scoreboard specialization(s)
//      Ex: typedef uvml_sb_simplex_c#(
//             .T_CNTXT(uvme_apb_timer_sb_cntxt_c),
//             .T_TRN  (uvma_apb_timer_mon_trn_c )
//          ) uvme_apb_timer_sb_simplex_c;

// Add tdefs, enums and structs here
// Ex: typedef bit [(`UVME_APB_TIMER_ABC_MAX_WIDTH-1):0]  uvme_apb_timer_abc_b_t;
// Ex: typedef enum {
//        UVME_APB_TIMER_MY_ABC
//     } uvme_apb_timer_my_enum;
// Ex: typedef struct {
//        bit [2:0]  abc;
//        logic      xyz;
//     } uvme_apb_timer_my_struct;


`endif // __UVME_APB_TIMER_TDEFS_SV__