// Copyright 2023 Acme Enterprises
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_CVMCU_IO_ST_BASE_TEST_WORKAROUNDS_SV__
`define __UVMT_CVMCU_IO_ST_BASE_TEST_WORKAROUNDS_SV__


// Temporary configuration constraints belong here (this file should be empty by the end of the project).


`endif // __UVMT_CVMCU_IO_ST_BASE_TEST_WORKAROUNDS_SV__