// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_CVMCU_IO_FTDECS_SV__
`define __UVMA_CVMCU_IO_FTDECS_SV__


typedef class uvma_cvmcu_io_cfg_c     ;
typedef class uvma_cvmcu_io_cntxt_c   ;
typedef class uvma_cvmcu_io_mon_trn_c ;
typedef class uvma_cvmcu_io_seq_item_c;
typedef class uvma_cvmcu_io_padi_mon_trn_c;
typedef class uvma_cvmcu_io_board_padi_seq_item_c;
typedef class uvma_cvmcu_io_chip_padi_seq_item_c;typedef class uvma_cvmcu_io_pado_mon_trn_c;
typedef class uvma_cvmcu_io_chip_pado_seq_item_c;
typedef class uvma_cvmcu_io_board_pado_seq_item_c;
typedef class uvma_cvmcu_io_mon_vseq_c ;
typedef class uvma_cvmcu_io_idle_vseq_c;
typedef class uvma_cvmcu_io_board_drv_vseq_c;
typedef class uvma_cvmcu_io_chip_drv_vseq_c;


`endif // __UVMA_CVMCU_IO_FTDECS_SV__