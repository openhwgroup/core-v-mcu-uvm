// Copyright 2022 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_UDMA_RX_DP_IN_TDEFS_SV__
`define __UVMA_UDMA_RX_DP_IN_TDEFS_SV__


// Add enums and structs here
// Ex: typedef bit [(`UVMA_UDMA_RX_DP_IN_ABC_MAX_WIDTH-1):0]  uvma_udma_rx_dp_in_abc_b_t;
// Ex: typedef enum {
//        UVMA_UDMA_RX_DP_IN_MY_ABC
//     } uvma_udma_rx_dp_in_my_enum;
// Ex: typedef struct {
//        bit [2:0]  abc;
//        logic      xyz;
//     } uvma_udma_rx_dp_in_my_struct;


`endif // __UVMA_UDMA_RX_DP_IN_TDEFS_SV__
