// Copyright 2024 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_APB_TIMER_SS_FTDECS_SV__
`define __UVMT_APB_TIMER_SS_FTDECS_SV__


`endif // __UVMT_APB_TIMER_SS_FTDECS_SV__