// Copyright 2023 Datum Technology Corporation
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_TCOUNTER_B_IF_CHKR_SV__
`define __UVMA_TCOUNTER_B_IF_CHKR_SV__


/**
 * Module encapsulating assertions targeting Timer unit counter Block Agent interface.
 * @ingroup uvma_tcounter_b_pkg
 */
module uvma_tcounter_b_if_chkr (
   uvma_tcounter_b_if  agent_if ///< Target interface
);

   // TODO Add assertions and/or functional coverage to uvme_tcounter_b_chkr

endmodule : uvma_tcounter_b_if_chkr


`endif // __UVMA_TCOUNTER_B_IF_CHKR_SV__