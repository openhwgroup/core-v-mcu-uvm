// Copyright 2023 Acme Enterprises
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_TPRESCALER_B_MACROS_SVH__
`define __UVMT_TPRESCALER_B_MACROS_SVH__


// Add preprocessor macros here
// Ex: `ifndef UVMT_TPRESCALER_B_ABC_WIDTH
//        `define UVMT_TPRESCALER_B_ABC_WIDTH 32
//     `endif


`endif // __UVMT_TPRESCALER_B_MACROS_SVH__