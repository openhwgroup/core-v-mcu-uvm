// Copyright 2022 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_UDMA_RX_MACROS_SVH__
`define __UVME_UDMA_RX_MACROS_SVH__


// Add preprocessor macros here
// Ex: `ifndef UVME_UDMA_RX_ABC
//        `define UVME_UDMA_RX_ABC 32
//     `endif


`endif // __UVME_UDMA_RX_MACROS_SVH__
