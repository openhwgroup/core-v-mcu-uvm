// Copyright 2023 Acme Enterprises
// All rights reserved.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMA_ADV_TIMER_B_CONSTANTS_SV__
`define __UVMA_ADV_TIMER_B_CONSTANTS_SV__


const int unsigned  uvma_adv_timer_b_default_num_bits  = 16; ///< Default  width.  Measured in bits (b).
const int unsigned  uvma_adv_timer_b_default_n_extsig  = 32; ///< Default  width.  Measured in bits (b).


`endif // __UVMA_ADV_TIMER_B_CONSTANTS_SV__